library ieee;
use ieee.std_logic_1164.all;

entity clkDiv is
	port(
		clk	: in std_ulogic;
		rst	: in std_ulogic;
		half_period : in std_ulogic;
		clk_out	: out std_ulogic
	);
end entity;

architecture clkDiv_arch of clkDiv is

	begin



end architecture;